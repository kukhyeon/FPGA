`timescale 1ns / 1ps
module mux_16to1v2(
    input   [3:0]   A,      // �Է� A (4��Ʈ)
    input   [3:0]   B,      // �Է� B (4��Ʈ)
    input   [3:0]   C,      // �Է� C (4��Ʈ)
    input   [3:0]   D,      // �Է� D (4��Ʈ)
    input   [3:0]   sel,    // ���� ��ȣ (4��Ʈ)
    output          Y       // ��� Y
    );
    
    wire out_8to1_1, out_8to1_2; // 8:1 ��Ƽ�÷��� ��� ��ȣ ����

    // ù ��° 8:1 ��Ƽ�÷��� �ν��Ͻ�
    mux_8to1 mux_8to1_1 (
        .a(A[1:0]),      // A�� ���� 2��Ʈ
        .b(A[3:2]),      // A�� ���� 2��Ʈ
        .c(B[1:0]),      // B�� ���� 2��Ʈ
        .d(B[3:2]),      // B�� ���� 2��Ʈ
        .sel(sel[2:0]),  // ���� 3��Ʈ ���� ��ȣ
        .out(out_8to1_1) // ù ��° 8:1 MUX ���
    );

    // �� ��° 8:1 ��Ƽ�÷��� �ν��Ͻ�
    mux_8to1 mux_8to1_2 (
        .a(C[1:0]),      // C�� ���� 2��Ʈ
        .b(C[3:2]),      // C�� ���� 2��Ʈ
        .c(D[1:0]),      // D�� ���� 2��Ʈ
        .d(D[3:2]),      // D�� ���� 2��Ʈ
        .sel(sel[2:0]),  // ���� 3��Ʈ ���� ��ȣ
        .out(out_8to1_2) // �� ��° 8:1 MUX ���
    );

    // ���� ��� ����: sel[3] ��Ʈ�� ���� �� 8:1 MUX �� �ϳ��� ����
    assign Y = (sel[3] == 0) ? out_8to1_1 : out_8to1_2;
endmodule
